module test(
    input [3:0]A,
    input [3:0]B,
    output reg [7:0]P
);




endmodule